-- IM : Instruction Memory --

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

entity IM is
    port(
        CLK : in std_logic;
        IMA : in std_logic_vector(31 downto 0);
        IMOut : out std_logic_vector(31 downto 0)
    );
end IM;

architecture RTL of IM is

begin
                  -- R Type : < op ><rs ><rt ><rd ><sha><func>
                  -- I Type : < op ><rs ><rt ><   imm/addr   >
                  -- J Type : < op ><          addr          >
    IMo : process(IMA(7 downto 2))
    begin
        case (IMA(7 downto 2)) is
        -- main:
            when "000000" =>  -- addi(1) rt(29),rs(29),-4
                    IMOut <= "000001"&"11101"&"11101"&"1111111111111100"; --4   --0
            when "000001" =>  -- sw(3) rt(31),rs(29),0
                    IMOut <= "000011"&"11101"&"11111"&"0000000000000000"; --8   --4
            when "000010" =>  -- addi(1) rt(3),rs(0),3
                    IMOut <= "000001"&"00000"&"00011"&"0000000000000011"; --04  --8
            when "000011" =>  -- jal(6) fact
                    IMOut <= "000110"&"00000000000000000000001000";       --18  --C
            when "000100" =>  -- sw(3),rt(2),rs(8),0
                    IMOut <= "000011"&"01000"&"00010"&"0000000000000000";  --0d  --10
            when "000101" =>  -- lw(2) rt(31),rs(29),0
                    IMOut <= "000010"&"11101"&"11111"&"0000000000000000";  --0b  --14
            when "000110" =>  -- addi(1) rt(29),rs(29),4
                    IMOut <= "000001"&"11101"&"11101"&"0000000000000100";  --07   --18
            when "000111" =>  -- jr(7) rs(31)
                    IMOut <= "000111"&"11111"&"000000000000000000000";      --1f  --1C
        -- fact:
            when "001000" =>  -- beq(4) rs(3),rt(0),return
                    IMOut <= "000100"&"00011"&"00000"&"0000000000001010"; --10  --20
            when "001001" =>  -- j(5) next
                    IMOut <= "000101"&"00000000000000000000001100";       --14  --24
        -- return:
            when "001010" =>  -- addi(1) rt(2),rs(0),1
                    IMOut <= "000001"&"00000"&"00010"&"0000000000000001"; 
            when "001011" =>  -- jr(7) rs(31)
                    IMOut <= "000111"&"11111"&"000000000000000000000";
        -- next
            when "001100" =>  -- addi(1) rt(29),rs(29),-8
                    IMOut <= "000001"&"11101"&"11101"&"1111111111111000"; --07  -30
            when "001101" =>  -- sw(3) rt(31),rs(29),4
                    IMOut <= "000011"&"11101"&"11111"&"0000000000000100"; --0F  --34
            when "001110" =>  -- sw(3) rt(3),rs(29),0
                    IMOut <= "000011"&"11101"&"00011"&"0000000000000000"; --0F  --38
            when "001111" =>  -- addi(1) rt(3),rs(3),-1
                    IMOut <= "000001"&"00011"&"00011"&"1111111111111111"; --04  --3C
            when "010000" =>  -- jal(6) fact
                    IMOut <= "000110"&"00000000000000000000001000";    --18 --40
            when "010001" =>  -- lw(2) rt(31),rs(29),4
                    IMOut <= "000010"&"11101"&"11111"&"0000000000000100"; --0b --44
            when "010010" =>  -- lw(2) rt(3),rs(29),0
                    IMOut <= "000010"&"11101"&"00011"&"0000000000000000"; --0b --48
            when "010011" =>  -- addi(1) rt(29),rs(29),8
                    IMOut <= "000001"&"11101"&"11101"&"0000000000001000"; --07 --4c
            when "010100" =>  -- mul rd(2),rs(3),rt(2)
                    IMOut <= "001000"&"00011"&"00010"&"00010"&"00000000000"; --20 --50
            when "010101" =>  -- jr(7) rs(31)
                    IMOut <= "000111"&"11111"&"000000000000000000000";        --1f  --54
            when others =>  -- nop : add $0,$0,$0
                    IMOut <= "00000000000000000000000000000000";
        end case;
    end process;

end RTL;